
module data_memory (clk,reset,we,addr,wd,rd);
input  clk, reset,we;
input



endmodule 